`timescale 1ns / 1ps

module PauseUnit(

	);
endmodule