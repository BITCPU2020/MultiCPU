`timescale 1ns / 1ps

module WRT(

    );
    
    mux #32 muxWD();
endmodule