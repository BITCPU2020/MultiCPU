`timescale 1ns / 1ps

module MultiCPU(

    );
    FTC ftc();
    DEC dec();
    EXE exe();
    MEM mem();
    WRT wrt();
endmodule