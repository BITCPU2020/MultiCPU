`timescale 1ns / 1ps

module MEM(

    ); 
    
    DataMemory data_memory();
    
endmodule
