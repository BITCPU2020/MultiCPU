`timescale 1ns / 1ps

module DataMemory(
		input wire clk, rstn,
		input wire i_DMem_dMemWe, i_DMem_sByte,
		input wire [31:0] i_DMem_addr,
		input wire [31:0] i_DMem_wData,
		output wire [31:0] o_DMem_rData
	);

	reg [7:0] dmem [255:0];

	// read
	wire [7:0] addr = i_DMem_addr[7:0];
	assign o_DMem_rData = (i_DMem_sByte == 1) ? {8'b0, 8'b0, 8'b0, dmem[addr]} :
						{dmem[addr+3], dmem[addr+2], dmem[addr+1], dmem[addr]};

	// write
	always @(posedge clk or negedge rstn) begin
		if (!rstn) begin
			dmem[0] <= 8'h0a;
			dmem[1]<=0;
			dmem[2]<=0;
			dmem[3]<=0;
			dmem[4]<=0;
			dmem[5]<=0;
			dmem[6]<=0;
			dmem[7]<=0;
			dmem[8]<=0;
			dmem[9]<=0;
			dmem[10]<=0;
			dmem[11]<=0;
			dmem[12]<=0;
			dmem[13]<=0;
			dmem[14]<=0;
			dmem[15]<=0;
			dmem[16]<=0;
			dmem[17]<=0;
			dmem[18]<=0;
			dmem[19]<=0;
			dmem[20]<=0;
			dmem[21]<=0;
			dmem[22]<=0;
			dmem[23]<=0;
			dmem[24]<=0;
			dmem[25]<=0;
			dmem[26]<=0;
			dmem[27]<=0;
			dmem[28]<=0;
			dmem[29]<=0;
			dmem[30]<=0;
			dmem[31]<=0;
			dmem[32]<=0;
			dmem[33]<=0;
			dmem[34]<=0;
			dmem[35]<=0;
			dmem[36]<=0;
			dmem[37]<=0;
			dmem[38]<=0;
			dmem[39]<=0;
			dmem[40]<=0;
			dmem[41]<=0;
			dmem[42]<=0;
			dmem[43]<=0;
			dmem[44]<=0;
			dmem[45]<=0;
			dmem[46]<=0;
			dmem[47]<=0;
			dmem[48]<=0;
			dmem[49]<=0;
			dmem[50]<=0;
			dmem[51]<=0;
			dmem[52]<=0;
			dmem[53]<=0;
			dmem[54]<=0;
			dmem[55]<=0;
			dmem[56]<=0;
			dmem[57]<=0;
			dmem[58]<=0;
			dmem[59]<=0;
			dmem[60]<=0;
			dmem[61]<=0;
			dmem[62]<=0;
			dmem[63]<=0;
			dmem[64]<=0;
			dmem[65]<=0;
			dmem[66]<=0;
			dmem[67]<=0;
			dmem[68]<=0;
			dmem[69]<=0;
			dmem[70]<=0;
			dmem[71]<=0;
			dmem[72]<=0;
			dmem[73]<=0;
			dmem[74]<=0;
			dmem[75]<=0;
			dmem[76]<=0;
			dmem[77]<=0;
			dmem[78]<=0;
			dmem[79]<=0;
			dmem[80]<=0;
			dmem[81]<=0;
			dmem[82]<=0;
			dmem[83]<=0;
			dmem[84]<=0;
			dmem[85]<=0;
			dmem[86]<=0;
			dmem[87]<=0;
			dmem[88]<=0;
			dmem[89]<=0;
			dmem[90]<=0;
			dmem[91]<=0;
			dmem[92]<=0;
			dmem[93]<=0;
			dmem[94]<=0;
			dmem[95]<=0;
			dmem[96]<=0;
			dmem[97]<=0;
			dmem[98]<=0;
			dmem[99]<=0;
			dmem[100]<=0;
			dmem[101]<=0;
			dmem[102]<=0;
			dmem[103]<=0;
			dmem[104]<=0;
			dmem[105]<=0;
			dmem[106]<=0;
			dmem[107]<=0;
			dmem[108]<=0;
			dmem[109]<=0;
			dmem[110]<=0;
			dmem[111]<=0;
			dmem[112]<=0;
			dmem[113]<=0;
			dmem[114]<=0;
			dmem[115]<=0;
			dmem[116]<=0;
			dmem[117]<=0;
			dmem[118]<=0;
			dmem[119]<=0;
			dmem[120]<=0;
			dmem[121]<=0;
			dmem[122]<=0;
			dmem[123]<=0;
			dmem[124]<=0;
			dmem[125]<=0;
			dmem[126]<=0;
			dmem[127]<=0;
			dmem[128]<=0;
			dmem[129]<=0;
			dmem[130]<=0;
			dmem[131]<=0;
			dmem[132]<=0;
			dmem[133]<=0;
			dmem[134]<=0;
			dmem[135]<=0;
			dmem[136]<=0;
			dmem[137]<=0;
			dmem[138]<=0;
			dmem[139]<=0;
			dmem[140]<=0;
			dmem[141]<=0;
			dmem[142]<=0;
			dmem[143]<=0;
			dmem[144]<=0;
			dmem[145]<=0;
			dmem[146]<=0;
			dmem[147]<=0;
			dmem[148]<=0;
			dmem[149]<=0;
			dmem[150]<=0;
			dmem[151]<=0;
			dmem[152]<=0;
			dmem[153]<=0;
			dmem[154]<=0;
			dmem[155]<=0;
			dmem[156]<=0;
			dmem[157]<=0;
			dmem[158]<=0;
			dmem[159]<=0;
			dmem[160]<=0;
			dmem[161]<=0;
			dmem[162]<=0;
			dmem[163]<=0;
			dmem[164]<=0;
			dmem[165]<=0;
			dmem[166]<=0;
			dmem[167]<=0;
			dmem[168]<=0;
			dmem[169]<=0;
			dmem[170]<=0;
			dmem[171]<=0;
			dmem[172]<=0;
			dmem[173]<=0;
			dmem[174]<=0;
			dmem[175]<=0;
			dmem[176]<=0;
			dmem[177]<=0;
			dmem[178]<=0;
			dmem[179]<=0;
			dmem[180]<=0;
			dmem[181]<=0;
			dmem[182]<=0;
			dmem[183]<=0;
			dmem[184]<=0;
			dmem[185]<=0;
			dmem[186]<=0;
			dmem[187]<=0;
			dmem[188]<=0;
			dmem[189]<=0;
			dmem[190]<=0;
			dmem[191]<=0;
			dmem[192]<=0;
			dmem[193]<=0;
			dmem[194]<=0;
			dmem[195]<=0;
			dmem[196]<=0;
			dmem[197]<=0;
			dmem[198]<=0;
			dmem[199]<=0;
			dmem[200]<=0;
			dmem[201]<=0;
			dmem[202]<=0;
			dmem[203]<=0;
			dmem[204]<=0;
			dmem[205]<=0;
			dmem[206]<=0;
			dmem[207]<=0;
			dmem[208]<=0;
			dmem[209]<=0;
			dmem[210]<=0;
			dmem[211]<=0;
			dmem[212]<=0;
			dmem[213]<=0;
			dmem[214]<=0;
			dmem[215]<=0;
			dmem[216]<=0;
			dmem[217]<=0;
			dmem[218]<=0;
			dmem[219]<=0;
			dmem[220]<=0;
			dmem[221]<=0;
			dmem[222]<=0;
			dmem[223]<=0;
			dmem[224]<=0;
			dmem[225]<=0;
			dmem[226]<=0;
			dmem[227]<=0;
			dmem[228]<=0;
			dmem[229]<=0;
			dmem[230]<=0;
			dmem[231]<=0;
			dmem[232]<=0;
			dmem[233]<=0;
			dmem[234]<=0;
			dmem[235]<=0;
			dmem[236]<=0;
			dmem[237]<=0;
			dmem[238]<=0;
			dmem[239]<=0;
			dmem[240]<=0;
			dmem[241]<=0;
			dmem[242]<=0;
			dmem[243]<=0;
			dmem[244]<=0;
			dmem[245]<=0;
			dmem[246]<=0;
			dmem[247]<=0;
			dmem[248]<=0;
			dmem[249]<=0;
			dmem[250]<=0;
			dmem[251]<=0;
			dmem[252]<=0;
			dmem[253]<=0;
			dmem[254]<=0;
		end else if(i_DMem_dMemWe) begin
			if(i_DMem_sByte==1) begin
				dmem[addr] <= i_DMem_wData[7:0];
				dmem[addr+1] <= dmem[addr+1];
				dmem[addr+2] <= dmem[addr+2];
				dmem[addr+3] <= dmem[addr+3];
			end else begin
				dmem[addr] <= i_DMem_wData[7:0];
				dmem[addr+1] <= i_DMem_wData[15:8];
				dmem[addr+2] <= i_DMem_wData[23:16];
				dmem[addr+3] <= i_DMem_wData[31:24];
			end
		end
	end
endmodule