`timescale 1ns / 1ps

module EXE(

    );
    ALU alu();
    mux #32 muxA1();
    mux #32 muxA2();
    mux #32 muxB();
endmodule
