`timescale 1ns / 1ps

module MultiCPU(

    );
    F f();
    DEC dec();
    EXE exe();
    MEM mem();
    WRT wrt();
endmodule
