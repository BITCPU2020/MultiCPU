`timescale 1ns / 1ps

module BranchUnit(

	);
endmodule