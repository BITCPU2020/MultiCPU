`timescale 1ns / 1ps

module F(

    );
    InstructionMemory instruction_memory();
    ProgramCounter program_counter();
endmodule
