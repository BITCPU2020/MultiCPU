`timescale 1ns / 1ps

module FTC(

    );
    InstructionMemory instruction_memory();
    ProgramCounter program_counter();
endmodule